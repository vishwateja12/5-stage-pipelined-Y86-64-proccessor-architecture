module F_RegisterBlock(clk,f_predPC,F_predPC);

input clk;

inout [63:0] f_predPC ;
output reg [63:0] F_predPC;




endmodule